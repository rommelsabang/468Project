module registerbank (en, R, q0, q1, q2, q3, q4, q5, q6, q7, q8, q9, q10, q11, q12, q13, q14, q15);
input [31:0] R;
input [15:0] en;
output reg [31:0] q0, q1, q2, q3, q4, q5, q6, q7, q8, q9, q10, q11, q12, q13, q14, q15;
always @*
begin
case (en)
16'b0000000000000001: q0 = R;
16'b0000000000000010: q1 = R;
16'b0000000000000100: q2 = R;
16'b0000000000001000: q3 = R;
16'b0000000000010000: q4 = R;
16'b0000000000100000: q5 = R;
16'b0000000001000000: q6 = R;
16'b0000000010000000: q7 = R;
16'b0000000100000000: q8 = R;
16'b0000001000000000: q9 = R;
16'b0000010000000000: q10 = R;
16'b0000100000000000: q11 = R;
16'b0001000000000000: q12 = R;
16'b0010000000000000: q13 = R;
16'b0100000000000000: q14 = R;
16'b1000000000000000: q15 = R;
endcase
end
endmodule