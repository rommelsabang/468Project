module register_bank(register,din,R0,R1,R2,R3,R4,R5,R6,R7,R8,R9,R10,R11,R12,R13,R14,R15);
input [15:0] register;
input [31:0] din;
output reg [31:0] R0,R1,R2,R3,R4,R5,R6,R7,R8,R9,R10,R11,R12,R13,R14,R15;

always@*
begin 

case(register)

16'b0000000000000001: R0=din;
16'b0000000000000010: R1=din;
16'b0000000000000100: R2=din;
16'b0000000000001000: R3=din;
16'b0000000000010000: R4=din;
16'b0000000000100000: R5=din;
16'b0000000001000000: R6=din;
16'b0000000010000000: R7=din;
16'b0000000100000000: R8=din;
16'b0000001000000000: R9=din;
16'b0000010000000000: R10=din;
16'b0000100000000000: R11=din;
16'b0001000000000000: R12=din;
16'b0010000000000000: R13=din;
16'b0100000000000000: R14=din;
16'b1000000000000000: R15=din;
endcase
end
endmodule

