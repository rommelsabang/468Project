module rr(num,in,out);
input [31:0] in;
input [4:0] num;
output reg[31:0] out;
always@*
begin
case (num)
5'b00001:out = {in[1-1:0],in[31:1]};
5'b00010:out = {in[2-1:0],in[31:2]};
5'b00011:out = {in[3-1:0],in[31:3]};
5'b00100:out = {in[4-1:0],in[31:4]};
5'b00101:out = {in[5-1:0],in[31:5]};
5'b00110:out = {in[6-1:0],in[31:6]};
5'b00111:out = {in[7-1:0],in[31:7]};
5'b01000:out = {in[8-1:0],in[31:8]};
5'b01001:out = {in[9-1:0],in[31:9]};
5'b01010:out = {in[10-1:0],in[31:10]};
5'b01011:out = {in[11-1:0],in[31:11]};
5'b01100:out = {in[12-1:0],in[31:12]};
5'b01101:out = {in[13-1:0],in[31:13]};
5'b01110:out = {in[14-1:0],in[31:14]};
5'b01111:out = {in[15-1:0],in[31:15]};
5'b10000:out = {in[16-1:0],in[31:16]};
5'b10001:out = {in[17-1:0],in[31:17]};
5'b10010:out = {in[18-1:0],in[31:18]};
5'b10011:out = {in[19-1:0],in[31:19]};
5'b10100:out = {in[20-1:0],in[31:20]};
5'b10101:out = {in[21-1:0],in[31:21]};
5'b10110:out = {in[22-1:0],in[31:22]};
5'b10111:out = {in[23-1:0],in[31:23]};
5'b11000:out = {in[24-1:0],in[31:24]};
5'b11001:out = {in[25-1:0],in[31:25]};
5'b11010:out = {in[26-1:0],in[31:26]};
5'b11011:out = {in[27-1:0],in[31:27]};
5'b11100:out = {in[28-1:0],in[31:28]};
5'b11101:out = {in[29-1:0],in[31:29]};
5'b11110:out = {in[30-1:0],in[31:30]};
5'b11111:out = {in[31-1:0],in[31:31]};
default:out = in;
endcase
end
endmodule